

`default_nettype none

////////////////////////////


/*
  see,
    https://www.eevblog.com/forum/projects/multislope-design/75/
    https://www.eevblog.com/forum/metrology/diy-high-resolution-multi-slope-converter/450/
    https://patentimages.storage.googleapis.com/e2/ba/5a/ff3abe723b7230/US5200752.pdf

    https://www.eevblog.com/forum/metrology/selecting-an-op-amp-for-integrator/
    https://www.eevblog.com/forum/metrology/7-5digit-diy-voltmeter/
*/

// advantage of macros over localparam enum, is that they generate errors if not defined.
// disdvantage is that it is easy to forget the backtick


// consider use one-hot encoding?


`define STATE_RESET_START    0

`define STATE_RESET          2
`define STATE_SIG_SETTLE_START 3
`define STATE_SIG_SETTLE    4
`define STATE_SIG_START     5
`define STATE_FIX_POS_START 6
`define STATE_FIX_POS       7
`define STATE_VAR_START     8
`define STATE_VAR           9
`define STATE_FIX_NEG_START 10
`define STATE_FIX_NEG       11
`define STATE_VAR2_START    12
`define STATE_VAR2          14
`define STATE_RUNDOWN_START 15
`define STATE_RUNDOWN       16

`define STATE_PRERUNDOWN_START 19
`define STATE_PRERUNDOWN    18

`define STATE_FAST_BELOW_START 20
`define STATE_FAST_BELOW    21

`define STATE_FAST_ABOVE_START 22
`define STATE_FAST_ABOVE    23




`define REFMUX_NONE        2'b00
`define REFMUX_POS         2'b01
`define REFMUX_NEG         2'b10
`define REFMUX_BOTH        2'b11






module adc_modulation (


  input           clk,
  input           reset_n,



  // comparator input
  input           cmpr_val,

  // perhaps rename p_cc_aperture, p_cc_fix  etc.
  input [32-1:0]  p_clk_count_aperture,   // considuer rename ru_aperture  or just clk_count_runup
  input [24-1:0]  p_clk_count_reset,      // useful if running stand-alone,
  input [24-1:0]  p_clk_count_fix,
  inout [24-1:0]  p_clk_count_var,

  input           p_use_slow_rundown,
  input           p_use_fast_rundown,
  input           p_active_sigmux,     // whether to swtich in the input signal


  // outputs
  output reg adc_measure_valid,           // indicate/assert completion, and valid measurement

  // now a wire
  output wire [ 8-1:0]  monitor,

  output reg sigmux,
  output reg rstmux,
  output reg [ 2-1:0]  refmux,            // reference current mux


  // TODO need better name. hi = disable comparator and enable latch
  // corresponds to hardware.
  output reg      cmpr_latch_ctl,


  ///////////

  /*

    Feb. 2026. we could really simplify this
    by moving all these outside the adc.
    - and read/ update them

  */


  // counts
  output reg [24-1:0] clk_count_rstmux,
  output reg [32-1:0] clk_count_refmux_neg,
  output reg [32-1:0] clk_count_refmux_pos,
  output reg [24-1:0] clk_count_refmux_both,
  output reg [32-1:0] clk_count_sigmux,
  output reg [32-1:0] clk_count_aperture,


  // stats
  output reg [24-1:0] stat_count_refmux_pos_up,
  output reg [24-1:0] stat_count_refmux_neg_up,
  output reg [24-1:0] stat_count_cmpr_cross_up,

  // nore
  output reg [24-1:0] stat_count_var_up,
  output reg [24-1:0] stat_count_var_down,
  output reg [24-1:0] stat_count_fix_up,
  output reg [24-1:0] stat_count_fix_down,
  output reg [24-1:0] stat_count_flip


);


  reg [5-1:0]   state = 0; // RESET_START;


  //////////////////////////////////////////////////////
  // counters and settings  ...

  reg [31:0]  clk_count_down;



  /////////////////////////


  // better name.  aperture_ok perhaps.
  reg in_runup;


  reg [2-1:0] cmpr_crossr;              // perhaps add _transition? or cmpr_

  wire cmpr_cross_up     = cmpr_crossr == 2'b10;
  wire cmpr_cross_down   = cmpr_crossr == 2'b01;
  wire cmpr_cross_any    = cmpr_cross_up || cmpr_cross_down ;



  reg [2-1:0] refmux_pos_cross;
  reg [2-1:0] refmux_neg_cross;

  wire refmux_pos_cross_up  = refmux_pos_cross == 2'b01;
  wire refmux_neg_cross_up  = refmux_neg_cross == 2'b01;




  assign monitor[0] = reset_n;
  assign monitor[1] = adc_measure_valid;

  // assign monitor[2] = sigmux;
  assign monitor[2] = in_runup;
  assign monitor[3] = (state == `STATE_FAST_ABOVE_START);
  assign monitor[4] = (state == `STATE_FAST_BELOW_START);
  assign monitor[5] = (state == `STATE_RUNDOWN);

  assign monitor[6] = 1'b0;
  assign monitor[7] = 1'b0;





  /*
      nov 12. 2023.
    we double flop.  for meta-stability.
    ie. avoid read/use twice in same block, and can be evaluated differently.
    perhaps review.
  */
  reg cmpr_val_last;

  always @(posedge clk)


    begin

      clk_count_down <= clk_count_down - 1;


      /* TODO nov 12. 2023.
        review why we do this. double flopping for stability on the clock edge.
        shouldn't matter?
      */
      // sample/bind comparator val once on clock edge. improves speed.
      cmpr_val_last <=  cmpr_val;


      cmpr_crossr               <= {cmpr_crossr[0], cmpr_val};

      // TODO change name ref_sw_pos_cross
      // instrumentation for switch transitions for both pos,neg (and both).
      refmux_pos_cross          <= { refmux_pos_cross[0], refmux[0] }; // old, new
      refmux_neg_cross          <= { refmux_neg_cross[0], refmux[1] };

      // TODO count_pos_trans or cross pos_  or just count_pos_trans
      // TODO must rename. actually represents count of each on switch transiton = count_ref_pos_on and count_ref_neg_on.
      if(refmux_pos_cross_up)
        stat_count_refmux_pos_up     <= stat_count_refmux_pos_up + 1;

      if(refmux_neg_cross_up)
        stat_count_refmux_neg_up     <= stat_count_refmux_neg_up + 1;

      if(cmpr_cross_up)
        stat_count_cmpr_cross_up     <= stat_count_cmpr_cross_up + 1;


      /*
        EI. use strategy of reading and counting the mux state values across the fsm state.
        avoids having to track for each state.
        ----
        it might also be more cycle accurate - given the phase transition setup, and comparator reads etc.
        but would need 32 bit values.
        - reduces spi overhead. if supported 32 byte reads.
        - reduces littering of count_var_up/count_var_down
        - reduces having to multiply out clk_count_var * count_var_up etc.
        - enables having non standar variable periods. eg. to reduce extra cycling to get to the other side.
        ------
            the way to evaluate is to use stderr(regression).
      */

      // synchronous behavior for all states

      case (refmux)

        `REFMUX_NEG:
            clk_count_refmux_neg <= clk_count_refmux_neg + 1;

        `REFMUX_POS:
            clk_count_refmux_pos <=  clk_count_refmux_pos + 1;

        `REFMUX_BOTH:
            begin
              clk_count_refmux_both <= clk_count_refmux_both + 1;
              clk_count_refmux_neg <= clk_count_refmux_neg + 1;
              clk_count_refmux_pos <=  clk_count_refmux_pos + 1;
            end

        `REFMUX_NONE:
          ; // switches are turned off at start. and also at prerundown.
            // don't really need to count this

      endcase



      if(rstmux)
        clk_count_rstmux <= clk_count_rstmux + 1;


      if(sigmux )
        clk_count_sigmux <= clk_count_sigmux + 1;


      if(in_runup)
        clk_count_aperture <= clk_count_aperture + 1;



      // runup termination condition
      if(clk_count_aperture >= p_clk_count_aperture)
        begin
          // stop signal input integration
          sigmux  <= 0;

          // indicate we finished RU
          in_runup <= 0;
        end



      ///////////////////////////////////

      case (state)


        `STATE_RESET_START:

          // reset state
          begin

            // setup next state to advance to if reset_n not asserted
            state           <= `STATE_RESET;

            // indicate no valid measurement available
            adc_measure_valid <= 0;

            clk_count_rstmux <= 0;   // clear rst count here

            clk_count_down  <= p_clk_count_reset;


            // hold integrator in reset
            in_runup        <= 0;
            sigmux          <= 0;
            rstmux          <= 1;
            refmux          <= `REFMUX_NONE;

            cmpr_latch_ctl  <= 1; // disable comparator, enable latch
          end



        `STATE_RESET:    // let integrator reset.
            if(clk_count_down == 0)
              state <= `STATE_SIG_START;



        // turn on signal integration, turn off reset, begin two phase runup
        `STATE_SIG_START:
          begin
            state                 <= `STATE_FIX_POS_START;

            // start input integration
            in_runup              <= 1;                     // start runup
            sigmux                <= p_active_sigmux;    // turn on signal input
            rstmux                <= 0;                     // turn off reset
            refmux                <= `REFMUX_NONE;          // keep refmux off

            // clear counts
            clk_count_refmux_neg  <= 0;
            clk_count_refmux_pos  <= 0;
            clk_count_refmux_both   <= 0;
            clk_count_sigmux      <= 0;
            clk_count_aperture    <= 0;

            /////////////////////////////
            // consider do this at reset/ done state.
            // clear the stat counts
            stat_count_var_up      <= 0;
            stat_count_var_down    <= 0;
            stat_count_fix_up      <= 0;
            stat_count_fix_down    <= 0;
            stat_count_refmux_pos_up    <= 0;
            stat_count_refmux_neg_up  <= 0;
            stat_count_flip        <= 0;
            stat_count_cmpr_cross_up <= 0;
          end


        // cycle +-ref currents, with/or without signal
        `STATE_FIX_POS_START:
          begin
            state             <= `STATE_FIX_POS;
            clk_count_down    <= p_clk_count_fix;

            stat_count_fix_down    <= stat_count_fix_down + 1;
            refmux            <= `REFMUX_POS; // initial direction

            cmpr_latch_ctl  <= 0; // enable comparator, // JA correct. 0 means it is transparent.
                                  // MUST do here, after we have driven away from the zero-cross,  rather than state_sig_start.
                                  // to reduce/ chance of comparator output oscillation
                                  // nov 16 2023.. actually we shave oscillation at start.
                                  // which is preturbing signal.
          end

        `STATE_FIX_POS:
          if(clk_count_down == 0)
            state <= `STATE_VAR_START;



        // variable direction
        `STATE_VAR_START:
          begin
            state             <= `STATE_VAR;
            clk_count_down    <= p_clk_count_var;

            if( cmpr_val_last)   // test below the zero-cross
              begin
                refmux        <= `REFMUX_NEG;  // add negative ref. to drive up.
                stat_count_var_up  <= stat_count_var_up + 1;
              end
            else
              begin
                refmux        <= `REFMUX_POS;
                stat_count_var_down <= stat_count_var_down + 1;
              end
          end



        `STATE_VAR:
          if(clk_count_down == 0)
            state <= `STATE_FIX_NEG_START;


        `STATE_FIX_NEG_START:
          begin
            state         <= `STATE_FIX_NEG;
            clk_count_down    <= p_clk_count_fix;

            stat_count_fix_up  <= stat_count_fix_up + 1;
            refmux        <= `REFMUX_NEG;
          end


        `STATE_FIX_NEG:
          // TODO add switch here for 3 phase modulation variation.
          if(clk_count_down == 0)
            state <= `STATE_VAR2_START;


        // variable direction
        `STATE_VAR2_START:
          ///////////
          // EXTR.  actually since we stopped injecting signal - it doesn't matter how many cycles we use to get above zero-cross.
          // and it will happen reasonably quickly. because of the bias.
          // so just keep running complete 4 phase cycles until we get a cross. rather than force positive vars.
          //////////
          begin
            state             <= `STATE_VAR2;
            clk_count_down    <= p_clk_count_var;

            if( cmpr_val_last) // below zero-cross
              begin
                refmux        <= `REFMUX_NEG;
                stat_count_var_up  <= stat_count_var_up + 1;
              end
            else
              begin
                refmux        <= `REFMUX_POS;
                stat_count_var_down <= stat_count_var_down + 1;
              end
          end

        /*
          E. IMPORTANT
          - solution to jump immediately to pre/rundown. without extra cycling.
            is just to keep adding up fix periods until above cross.

        */
        `STATE_VAR2:
          if(clk_count_down == 0)
            begin
              // runup already finished.
              if( !in_runup)

                if(p_use_fast_rundown)
                  begin
                    if(  cmpr_val_last) // below cross
                      state <= `STATE_FAST_BELOW_START;
                    else                      // above cross
                      state <= `STATE_FAST_ABOVE_START;
                  end
                else
                  begin
                    // above cross and last var was up phase
                    /*
                      TODO fixme. nov  2023. state removed.
                    */
                    if( refmux  == `REFMUX_NEG && ! cmpr_val_last)
                      state <= `STATE_PRERUNDOWN_START;
                    else
                      // keep cycling
                      state <= `STATE_FIX_POS_START;

                      stat_count_flip <= stat_count_flip + 1;
                  end

              // signal integration not finished
              else
                  // do another cycle
                  state <= `STATE_FIX_POS_START;
            end

        //////////////////////////////////////////////
        // fast rundown.

        /*
        EXTR. cmpr hysteresis. affects setup for rundown.
        means we don't have to pad small extra clk count,
        to guarantee, we don't miss a crossing.
        */
        // we are somewhere above zero,
        // advance until below zero cross.
        `STATE_FAST_ABOVE_START:
          begin
            refmux          <= `REFMUX_POS;

            if( cmpr_val_last)                  // below zero-cross. EXTR. note not a comparator transition test. instead an actual value .
              state   <= `STATE_FAST_BELOW_START;     // advance to below_start.
          end


        /*
          cmpr hystersis means more clk cycles, than  would need for exact cross.
          also slope-amp will determine how many clk cycles needed to get across positive hysterisis.

        */
        // advance until above zero-cross.
        `STATE_FAST_BELOW_START:
           begin
            refmux    <= `REFMUX_NEG;

             if( ! cmpr_val_last) // above zero-cross
              begin
                state         <= `STATE_RUNDOWN_START; // goto rundown.

                /* nov 20, 2023.
                  turn off both +ve and -ve currents, to equalize switch counts and charge-injection - for +ve and -ve ref.
                - This code should be kept. because a half-wave switch has far more charge-injection - that full-wave on/off cycle - where most will be cancelled.
                  and this applies - if the sequence is spread over two switches - for both +ref and -ref currents..
                  reduces noise.  0.7uV to 0.6uV or lower. RMS 1nplc .
                --
                - remember abrupt chages in noise, are due to variations in run-up counts, between measurements due to slight thermal shifts.
                */
                refmux    <= `REFMUX_NONE;
              end
            end






        `STATE_RUNDOWN_START:
          begin
            state         <= `STATE_RUNDOWN;

            /*
              IMPORTANT. we are not counting a possible switch transition here.
              Bug?
            */
            if( p_use_slow_rundown )
              // turn on both references - to create +ve bias, to drive integrator down.
              refmux      <= `REFMUX_BOTH;
            else
              // fast rundown
              refmux      <= `REFMUX_POS;
          end


        `STATE_RUNDOWN:
          begin
            // TODO change to cmpr_val test.
            // zero-cross to finish. should probably change to use last_comparator
              /*
              EXTR. at rundown, even though we approach from same direction,
              we may get a cross in either direction (up/down) due to cmpr glitching.
              this applies even if usign the cmpr latch, because the latch only guarantees hold, not value, and has a delay
              So must check in both directions.
              hysterisis works as a practical solution
              --
              - using external ff to control cmpr latch, may even hide a transition from being seen by fpga. so is not a solution.
              - unless use the ff output.
              */

            if(cmpr_cross_any )
              begin

                cmpr_latch_ctl          <= 1; // disable comparator,

                // signal valid measurement.
                adc_measure_valid <= 1;

                // next transition
                state                   <= `STATE_RESET_START;


                // hold in reset
                in_runup        <= 0;
                sigmux          <= 0;
                rstmux          <= 1;
                refmux          <= `REFMUX_NONE;

/*
                // counts
                clk_count_rstmux_last       <= clk_count_rstmux;    // this doesn't work. reports 0.
                clk_count_refmux_neg_last   <= clk_count_refmux_neg;
                clk_count_refmux_pos_last   <= clk_count_refmux_pos;
                clk_count_refmux_both_last  <= clk_count_refmux_both;
                clk_count_sigmux_last       <= clk_count_sigmux;
                clk_count_aperture_last     <= clk_count_aperture;

                // stats
                stat_count_refmux_pos_up_last <= stat_count_refmux_pos_up;
                stat_count_refmux_neg_up_last <= stat_count_refmux_neg_up;
                stat_count_cmpr_cross_up_last <= stat_count_cmpr_cross_up;

                stat_count_var_up_last      <= stat_count_var_up;
                stat_count_var_down_last    <= stat_count_var_down;
                stat_count_fix_up_last      <= stat_count_fix_up;
                stat_count_fix_down_last    <= stat_count_fix_down;
                stat_count_flip_last        <= stat_count_flip;
*/

                // stat_clk_count_rundown_last  <= clk_count;                           // why do we record this

              end
          end

      endcase



      // override all states - if reset_n enabled, then don't advance out-of reset state.
      if(reset_n == 0)      // in reset
        begin

            state <= 0;
        end



    end


endmodule


