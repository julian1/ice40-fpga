
/*
  - can have heartbeat timer. over spi.
      but don't want to spew spi tranmsission during acquisition.

  - if have more than one dac. then just create another register. very clean.
   - perhaps instead of !cs or !cs2.  could write macro  or asserted_n(cs ) etc
*/



// `include "../../common/mux_spi.v"
`include "../../common/mux_assign.v"
`include "../../common/test_pattern.v"
`include "../../common/timed_latch.v"

`include "register_set.v"
`include "sample_acquisition_pc.v"

`include "sample_acquisition_az.v"

`include "adc-mock.v"       // change name adc-mock.
`include "refmux-test.v"

`include "adc_modulation_05.v"
`include "sample_acquisition_no_az.v"
`include "sequence_acquisition.v"

`default_nettype none



module top (

  // these are all treated as wires.

  // input  CLK,


  ////////////////////////
  // spi

  /*#A dual-function, serial output pin in both configuration modes.
  #iCE40 LM devices have this pin shared with hardened SPI IP
  #SPI_MISO pin. */
  output SDO,

  /*# A dual-function, serial input pin in both configuration modes.
  # iCE40 LM devices have this pin shared with hardened SPI IP
  # SPI_MOSI pin. */
  input SDI,

  /*#A dual-function clock signal. An output in Master mode and
  #input in Slave mode. iCE40 LM devices have this pin shared with
  # hardened SPI IP SPI_SCK pin.*/
  input SCK,

  /*#An important dual-function, active-low slave select pin. After
  #the device exits POR or CRESET_B is toggled (High-Low-High), it
  #samples the SPI_SS to select the configuration mode (an output
  #in Master mode and an input in Slave mode). iCE40 LM devices
  #have this pin shared with hardened SPI IP SPI1_CSN pin.*/
  input SS,


  input  SPI_CS2,


  ///////////
  output [ 4-1: 0 ] leds_o,

  output [ 8-1: 0]  monitor_o,

  input [4-1: 0]    hw_flags_i,



  input  CLK,




  // 4094
  output GLB_SPI_MOSI,
  output GLB_SPI_CLK,
  output GLB_4094_OE_CTL,
  output GLB_4094_STROBE_CTL,

  output SPI_DAC_SS,

  input U1004_4094_DATA,


  input trigger_source_external_i,   // trigger_ext_out   - need to re
  input trigger_source_internal_i,   // trigger_int_out 38
  input unused1_i,                    // 39


  output spi_interrupt_ctl_o,
  output meas_complete_o,


  // output sig_pc1_sw_o,
  // output sig_pc2_sw_o ,

  output [ 2-1: 0 ] pc_sw_o,

  // az mux
  // u410
  output [ 4-1: 0 ] azmux_o,


  // adc comparator latch ctl.
  // should be cmpr_latch_ctl
  output adc_cmpr_latch_ctl_o,

  input adc_cmpr_p_i,


  // U902. adc ref current mux
  output [ 4-1: 0 ] adc_refmux_o,

/*


  //
  // inputs

  // spi
  input  SPI_CLK,
  input  SPI_CS,
  input  SPI_MOSI,
  input  SPI_CS2,
  output SPI_MISO,
  // output b

  input U1004_4094_DATA,
  input LINE_SENSE_OUT,
  input SWITCH_SENSE_OUT,
  input DCV_OVP_OUT,
  input OHMS_OVP_OUT,
  input SUPPLY_SENSE_OUT,
  input UNUSED_2,                    // change name UNUSED_2_OUT

  // input  U1004_4094_DATA,   // this is unused. but it's an input


  //
  output SPI_INTERRUPT_CTL,    // should be modeal. eg. same as meas complete
  output MEAS_COMPLETE_CTL,

  //  adc current switches
  output U902_SW0_CTL,
  output U902_SW1_CTL,
  output U902_SW2_CTL,
  output U902_SW3_CTL,
  output CMPR_LATCH_CTL,

  ////////////
*/

);




  ////////////////////////////////////////
  // spi muxing

  /*
    TODO. rather than pulling all these out in vectors.
          we should combine in line/place. the same way we do mux align.
          eg.

      . vec_cs(  {  dummy,  GLB_4094_STROBE_CTL  }   ),
      ote. we are already doing this for polarity
  */

  wire [32-1:0] reg_spi_mux ;// = 8'b00000001; // test

  assign GLB_SPI_CLK          = reg_spi_mux == 8'b0 ? 1 : SCK;      // park hi

  assign GLB_SPI_MOSI         = reg_spi_mux == 8'b0 ? 1 : SDI;      // park hi

  assign GLB_4094_STROBE_CTL  = reg_spi_mux == 8'b01 ?  (~ SPI_CS2)  : 0;     // active hi

  assign SPI_DAC_SS           = reg_spi_mux == 8'b10 ?  SPI_CS2 : 1;     // active lo


  wire w_dout ;

  assign w_dout = SDO;




/*
  // would be nice to project these in a mode,
  // but if there's a spi problem - we are unlikely to get it into a mode.

  assign monitor_o[0]  = GLB_SPI_CLK;
  assign monitor_o[1]  = GLB_SPI_MOSI;
  assign monitor_o[2]  = SPI_DAC_SS     ;
*/




  /////////////////////////////////////////////
  // 4094 OE
  wire [32-1:0] reg_4094;   // TODO rename
  assign { GLB_4094_OE_CTL } = reg_4094;    //  lo. start up not enabled.

  ////////////////////////////////////////



  wire [32-1:0] reg_direct;

  // wire [32-1 :0] reg_sa_arm_trigger;              // only a single bit is needed here. should be able to write to handle more efficiently.




  // readable inputs
  wire [32 - 1 :0] reg_status ;

  assign reg_status = {



    21'b0,

    hw_flags_i,

    { 8'b10101010 }  // magic
/*
    8'b0 ,
    monitor,                          // don't see having the monitor readable through a different register is useful.   a git commit or crc would be useful.
                                      // add a count, as a transactional read lock.
    HW2,  HW1,  HW0,

    reg_sa_arm_trigger[0],            // ease having to do a separate register read, to retrieve state.
    sample_acquisition_az_status_out, // 3 bits
    adc2_measure_valid,

    // HW2,  HW1,  HW0 ,   4'b0,  outputs_vec[ `IDX_SPI_INTERRUPT_CTL ] ,

    3'b0,
    SWITCH_SENSE_OUT, DCV_OVP_OUT, OHMS_OVP_OUT, SUPPLY_SENSE_OUT, UNUSED_2
*/
 };


  // verilog literals are hard!.
  // 4'b1                         == 0001
  // { 1,1,1,1}                   == 0001
  // { 1'b1, 1'b1, 1'b1, 1'b1 }   == 1111
  // 4 { 1'b1 }                   == 1111
  // 4'b1111                      == 1111

  wire [32-1 :0] reg_mode;     // _mode or AF reg_af alternate function  two bits




  // TODO drop the _out suffix. because any wire is a driver in the context of the top module.
  // should prefix o_test_pattern ?  or just on module names?
  wire [32-1 :0] test_pattern_out;

  test_pattern  test_pattern_1 (
    . clk( CLK),
    . out( test_pattern_out)
  );




  wire [32-1:0] reg_sa_p_clk_count_precharge;

  wire [32-1:0] reg_sa_p_seq_n;
  wire [32-1:0] reg_sa_p_seq0;
  wire [32-1:0] reg_sa_p_seq1;
  wire [32-1:0] reg_sa_p_seq2;
  wire [32-1:0] reg_sa_p_seq3;


  wire [32-1 :0] reg_adc_p_clk_count_aperture;  // 32/31 bit nice. for long sample.
  wire [32-1 :0] reg_adc_p_clk_count_reset;

  ////////
  // rename sa_simple_ ?
  // sa_pc_test
  // or test_sa_pc

  /*
    - note that we can still hook this up to the adc. for measurement.
    - slightly different from a direct mode. where there is no pc switching.

    TODO. rename include test in name. it's actually sample acquisition.
  */


/*
      ================
    - EXTR.  NOT clear we even need the sample_acquisition_pc   - because can just use the sequence-acquisition.
          and keep the azmux held off.
        or even the non mocked.
      eg.  i think the sample sequence controller - can manage to encode the pc  switching test.  also. by just holding the azmux off.
    ================
*/

  wire sample_acquisition_pc_sw_pc_ctl;
  wire sample_acquisition_pc_led0;
  wire [8-1 : 0] sample_acquisition_pc_monitor;


  // rename this doesn't do sample acquisition. it just switches the pre-charge
  // we will switch to another mode  - before and after - in order to measure charge contribution

  sample_acquisition_pc
  sample_acquisition_pc (
    // inputs
    .clk(CLK),
    .reset_n( 1'b0 ),                       // JA. EXTR. consider placing the bit in output reg. so that it can be enabled in the corresponding mode.
                                            // likewise should be able to activate the adc in direct mode, by flipping the bit.  except won't work. because doesn't have control over refmux, comparator etc.
                                            // But may be useful to create a direct mode (with no sequence), but with the adc.
                                            // ---
                                            // or connect to the trigger. because the behavior is much the same - as the sequence controller.

    // inputs
    .p_clk_sample_duration_i( reg_adc_p_clk_count_aperture ),
    .p_clk_count_precharge_i( reg_sa_p_clk_count_precharge[ 24-1:0] ),

    // outputs
    .sw_pc_ctl_o( sample_acquisition_pc_sw_pc_ctl   ),          // should pass in both. and a register like a mask. to indicate which to use. similar to register for az mux.  might encode in same register.
    .led0_o(      sample_acquisition_pc_led0 ),                 // EXTR. just use the bits of reg_direct for azmux and which pc switch to use.  add back reg_direc2 for the ratiometric.
    .monitor_o(   sample_acquisition_pc_monitor  )
  );






  ////////////////////////

  wire          adc_mock_reset_n;
  wire          adc_mock_measure_valid;
  wire [8-1:0 ] adc_mock_monitor;

  adc_mock
  adc_mock (

    .clk(CLK),
    .reset_n( adc_mock_reset_n ),

    // inputs
    .p_clk_count_aperture_i( reg_adc_p_clk_count_aperture ),

    // outputs
    .adc_measure_valid_o( adc_mock_measure_valid ),
    .monitor_o(  adc_mock_monitor )
  );


  // fucking hell it's getting a bit complicated.
  // we need to rename this.   sa_az_adc_mock_sw_pc_ctl.
  wire [2-1:0]  sample_acquisition_az_sw_pc_ctl;
  wire [4-1:0]  sample_acquisition_az_azmux;

  wire [4-1:0]  sample_acquisition_az_leds;
  wire [8-1:0]  sample_acquisition_az_monitor;
  wire [3-1:0]  sample_acquisition_az_status;
  // wire          sample_acquisition_az_adc_measure_trig;

/*
  sample_acquisition_az
  sample_acquisition_az (

    .clk(CLK),
    .reset_n( trigger_source_internal_i ),    // we want this to remove. the old edge triggered stuff.

    // inputs
    .adc_measure_valid_i( adc_mock_measure_valid ),                     // fan-in from adc

    // TODO move to registers
    .p_seq0_i( reg_sa_p_seq0[ 4-1:0]  ),
    .p_seq1_i( reg_sa_p_seq1[ 4-1:0]  ),
    .p_seq2_i( reg_sa_p_seq2[ 2-1:0] ),
    .p_clk_count_precharge_i( reg_sa_p_clk_count_precharge[ 24-1:0]  ),     // done

    // outputs
    .sw_pc_ctl_o( sample_acquisition_az_sw_pc_ctl  ),
    .azmux_o (    sample_acquisition_az_azmux  ),
    .led0_o(      sample_acquisition_az_led0  ),
    .monitor_o(   sample_acquisition_az_monitor  ),    // only pass 2 bit to the az monitor
    .status_o(  sample_acquisition_az_status ),

    .adc_reset_no(  adc_mock_reset_n  )
  );
*/

  // rename sample_acquisition_sequence
  sequence_acquisition
  sequence_acquisition (

    .clk(CLK),
    .reset_n( trigger_source_internal_i ),    // we want this to remove. the old edge triggered stuff.

    // inputs
    .adc_measure_valid_i( adc_mock_measure_valid ),                     // fan-in from adc


    // TODO move to registers

    .p_seq_n_i( reg_sa_p_seq_n[ 2-1: 0]  ),
    .p_seq0_i( reg_sa_p_seq0[ 6-1: 0]  ),
    .p_seq1_i( reg_sa_p_seq1[ 6-1: 0]  ),
    .p_seq2_i( reg_sa_p_seq2[ 6-1: 0] ),
    .p_seq3_i( reg_sa_p_seq2[ 6-1: 0] ),


    .p_clk_count_precharge_i( reg_sa_p_clk_count_precharge[ 24-1:0]  ),     // done

    // outputs
    .sw_pc_ctl_o( sample_acquisition_az_sw_pc_ctl  ),
    .azmux_o (    sample_acquisition_az_azmux  ),

    .leds_o(      sample_acquisition_az_leds  ),
    .monitor_o(   sample_acquisition_az_monitor  ),    // only pass 2 bit to the az monitor
    .status_o(  sample_acquisition_az_status ),

    .adc_reset_no(  adc_mock_reset_n  )
  );


  ////////////////////




















  /////////////////////////
  // We could do one led, for SS, and one for CS2 (4094,etc).
  // rename timed_latch_hold
  /*
    change name. this delay stretch the signal over longer clk duration.
  */
  wire led0;
  timed_latch timed_latch (
    . clk(CLK),
    . trig_i( !SS || !SPI_CS2 ),      // rename set?
    . out( led0 )
  );



  // TODO consider rename adc_refmux_test.
  wire [8-1:0] refmux_test_monitor;
  wire [4-1:0] refmux_test_refmux;

  refmux_test refmux_test (

    .clk(CLK),
    // JA.   add a reset_n.  and only activate in the corresponding mode.
    // we don't care about reset here

    . p_clk_count_reset_i( $rtoi(  `CLK_FREQ * 500e-6 )  ), // 500us.
    . p_clk_count_fix_i(   $rtoi( `CLK_FREQ * 100e-6 )) ,  // 100us. initial but too long

    . cmpr_val_i( adc_cmpr_p_i ),

    .monitor_o( refmux_test_monitor),
    /* ie. refmux order pos,neg,source,reset.
      do we want to change this in main.pcf.. no keep ic sw pinout order.  */
    .refmux_o ( { refmux_test_refmux[  3  ],  refmux_test_refmux[ 0 +: 2 ]   }  ),
    .sigmux_o( refmux_test_refmux[ 2] )
  );







  ////////////////////////////

  // adc gets instantiated once, so should be called adc. not adc2.
  // do the no_az first. as the simplest.

  // TODO rename adc
  wire          adc2_reset_n;
  wire          adc2_measure_valid;

  wire [8-1: 0 ] adc2_monitor;
  wire [4-1: 0 ] adc2_mux;
  wire           adc2_cmpr_latch_ctl;


  wire [24-1:0] adc2_clk_count_refmux_reset_last;
  wire [32-1:0] adc2_clk_count_refmux_neg_last;    // maybe add reg_ prefix. No. they are not registers, until they are in the register_bank context.
  wire [32-1:0] adc2_clk_count_refmux_pos_last;
  wire [24-1:0] adc2_clk_count_refmux_rd_last;
  wire [32-1:0] adc2_clk_count_mux_sig_last;

  wire [24-1 :0] adc2_stat_count_refmux_pos_up_last;
  wire [24-1 :0] adc2_stat_count_refmux_neg_up_last;
  wire [24-1 :0] adc2_stat_count_cmpr_cross_up_last;


  adc_modulation
  adc2(

    .clk(CLK),
    .reset_n( adc2_reset_n),      // OK.


    .cmpr_val( adc_cmpr_p_i ),                  // OK.  fan in-  rename top_adc_cmpr_p_i ?

    . p_clk_count_aperture( reg_adc_p_clk_count_aperture /*reg_adc_p_aperture */),
    . p_clk_count_reset( reg_adc_p_clk_count_reset[ 24-1: 0  ]  ) ,
    // . p_clk_count_fix( 24'd15 ) ,         // +-15V. reduced integrator swing.
    // . p_clk_count_var( 24'd100 ) ,

    . p_clk_count_fix( 24'd67 ) ,           // 1.5nF. 4x counts of 330p. oct. 2023. test.
    . p_clk_count_var( 24'd450 ) ,

    . p_use_slow_rundown( 1'b1 ),
    . p_use_fast_rundown( 1'b1 ),

    // outputs - ctrl
    .adc_measure_valid( adc2_measure_valid),    // OK, fan out back to the sa controllers
    .cmpr_latch_ctl( adc2_cmpr_latch_ctl   ),
    .monitor(  adc2_monitor  ),
    .refmux(  { adc2_mux[  3  ],  adc2_mux[ 0 +: 2 ]   } ),           // pos, neg, reset. are on two different 4053,
    .sigmux(    adc2_mux[  2  ] ),                                    // perhaps clearer if split into adcrefmux and adcsigmux in the wire assignment. but it would then need two vars.
                                                                      // which isn't representative of the single synchronizer. so do it here instead.
    // adc clk counts for last sample measurement
    .clk_count_refmux_reset_last(adc2_clk_count_refmux_reset_last),
    .clk_count_refmux_neg_last(  adc2_clk_count_refmux_neg_last),
    .clk_count_refmux_pos_last(  adc2_clk_count_refmux_pos_last),
    .clk_count_refmux_rd_last(   adc2_clk_count_refmux_rd_last),
    .clk_count_mux_sig_last(  adc2_clk_count_mux_sig_last ),

    // stats
    .stat_count_refmux_pos_up_last( adc2_stat_count_refmux_pos_up_last),
    .stat_count_refmux_neg_up_last( adc2_stat_count_refmux_neg_up_last),
    .stat_count_cmpr_cross_up_last( adc2_stat_count_cmpr_cross_up_last)
  );



  // wire [ `NUM_BITS-1:0 ]  sample_acquisition_no_az_out ;  // beter name ... _outputs_vec ?

  // wire sample_acquisition_no_az_reset_n;

  wire sample_acquisition_no_az_adc2_reset_n;
  wire sample_acquisition_no_az_led0 ;
  wire [8-1:0] sample_acquisition_no_az_monitor;


  // JA remove
  // new sequence controller should be able to handle,  by only sampling hi, with or without precharge switching, controlled with flags
  sample_acquisition_no_az
  sample_acquisition_no_az (

    .clk(CLK),
    .reset_n( trigger_source_internal_i ),

    // inputs
    .adc_measure_valid( adc2_measure_valid ),                     // fan-in from adc

    .p_clk_count_precharge( reg_sa_p_clk_count_precharge[ 24-1:0 ]),

    // outputs
    .led0(      sample_acquisition_no_az_led0  ),
    .monitor(   sample_acquisition_no_az_monitor  ),    // we could pass subset of monitor if watned. eg. only 4 pins...
    .adc_reset_no ( sample_acquisition_no_az_adc2_reset_n),
  );




  /*
      - It may be possible to control and run the adc - with the direct register. just be setting the bit for the trigger.
      - BUT. wants to be non edge triggered.

  */


  ////////////////////////////
  // unused. should be able to be wire?
  reg [32-26- 1:0] dummy_bits_o ;


  // mode, alternative function selection
  mux_8to1_assign #( 32  )
  mux_8to1_assign_1  (

    .a(  reg_direct  ),                         // mode/AF 0  MODE_DIRECT       note, could change to project the the spi signals on the monitor, for easier ddebuggin. no. because want direct to control all outputs for test.

    /* TODO remove.
        the modes for output lo, and output hi - are not really needed. eg. mode 0; direct 0xffffffff ; or 0x00000000; etc.
        and there maybe chance of damage, if parts are populated
      */
    .b(  32'b0  ),                              // mode/AF  1 MODE_LO           all outputs low.
    .c( { 32 { 1'b1 } }    ),                   // mode/AF 2  MODE_HI           all outputs hi.
    .d( test_pattern_out ),                     // mode/AF 3  MODE_PATTERN      pattern. needs xtal.

    // mode/AF 4 MODE_PC_TEST
    .e( {  { 32 - 14 { 'b0 }},
                                             // 14
          sample_acquisition_pc_sw_pc_ctl,  // 12+2
          sample_acquisition_pc_monitor,    // 4+8
          3'b0,                             // 1+3    - should be reg_direct.
          sample_acquisition_pc_led0        // 0+1
        } ),

/*
    .a( { 1'b0, { 15 { 1'b0 } },  reg_led[ 0], { 13 { 1'b0 } } }    ),        // 0. default mode. 0 on all outputs, except follow reg_led, for led.
    .b( { 1'b0, { `NUM_BITS { 1'b1 } } } ),             // 1.
    .c( { 1'b0, test_pattern_out } ),                   // 2
    .d( { 1'b0, reg_direct[ `NUM_BITS - 1 :  0 ]  } ), // 3.    // direct mode. register control.
    .e( { 1'b0, sample_acquisition_pc_out} ),                   // 4
    .f( { sample_acquisition_az_adc2_reset_n,    sample_acquisition_az_out } ),                   // 5
    .g( { sample_acquisition_no_az_adc2_reset_n, sample_acquisition_no_az_out } ),                // 6
    // .h( { 1'b0, { `NUM_BITS { 1'b1 } } } ),             // 7
    .h( { 1'b0, sa_no_az_test_out } ),             // 7
*/

    // mode/AF  5  MODE_AZ_TEST with a mocked adc.  useful. for timing/ control tests
    // very useful - allows testing precharge/az switching, even if don't have adc populated
    .f( {  { 32 - 26 { 'b0 }},
                                                // 26
          1'b0, // adc2_reset_n         // 25 + 1
          1'b0, // meas_complete              // 24+1
          1'b0,   // spi_interupt             // 23 + 1
          1'b0,  // adc_cmpr_latch            // 22+1
          4'b0,  // adc_refmux               // 18+4
          sample_acquisition_az_azmux,        // 14+4
          sample_acquisition_az_sw_pc_ctl,   // 12+2
          // adc_mock_monitor[0 +: 6] , sample_acquisition_az_monitor[ 0 +: 2],    // 4+8
          sample_acquisition_az_monitor[ 0 +: 8],    // 4+8
          sample_acquisition_az_leds        // 0+1
        } ),


    // mode  6. adc refmux test
    // limited modulation of ref currents, useful when populating pcb, don't need slope-amp/comparator etc.
    .g( {  { 32 - 22 { 'b0 }},
                                              // 22
          refmux_test_refmux,                // 18+4
          4'b0,    // azmux                  // 14+4
          2'b0 ,  // precharge               // 12+2
          refmux_test_monitor,            //     4+8
          4'b0   // leds                   // 0+4
        } ),


    // mode 7. full adc/ no az.
    .h( {  { 32 - 26 { 'b0 }},
                                                // 26
          sample_acquisition_no_az_adc2_reset_n,        // 25 + 1
          adc2_measure_valid,   // meas_complete              // 24+1
          adc2_measure_valid,   // spi_interupt   // 23 + 1
          adc2_cmpr_latch_ctl,  // adc_cmpr_latch   // 22+1
          adc2_mux,             // adc_refmux     // 18+4
          // use reg_direct to control the azmux
          reg_direct [ 14 +: 4 ],  // azmux      // 14+4
          2'b0 ,                  // precharge    // 12+2     // TODO fixme. samples boot only.  use reg_sa_p_pc.
          adc2_monitor[ 0 +: 6], sample_acquisition_no_az_monitor[ 0 +: 2],    // 4+8
          // 3'b0,                             // 1+3
          sample_acquisition_az_leds        // 0+1
        } ),



    .sel( reg_mode[ 3-1 : 0 ]),

    // leds and monitor go first, since they are the most generic functionality

    .out( {   dummy_bits_o,               // 26

              adc2_reset_n,        // 25 + 1

              meas_complete_o,          // 24+1     // interupt_ctl *IS* generic so should be at start, and connects straight to adum. so place at beginning. same argument for meas_complete
              spi_interrupt_ctl_o,      // 23+1     todo rename. drop the 'ctl'.
              adc_cmpr_latch_ctl_o,         // 22+1
              adc_refmux_o,             // 18+4     // better name adc_refmux   adc_cmpr_latch
              azmux_o,                  // 14+4
              pc_sw_o,              // 12+2
              monitor_o,                // 4+8
              leds_o                    // 0+4
            }  )

  );







  register_set // #( 32 )
  register_set
    (

    // should prefix fields with spi_
    . clk(   SCK ),
    . cs_n(  SS /*SPI_CS */ ),        // rename cs_n
    . din(   SDI /*SPI_MOSI */),


    . dout( w_dout ),            // drive miso from via muxer
    // . dout( SDO /* SPI_MISO */ ),        // drive miso output pin directly.


    // outputs
    . reg_spi_mux(reg_spi_mux),
    . reg_4094(reg_4094 ) ,
    . reg_mode(reg_mode),
    . reg_direct(reg_direct),

    // inputs
    . reg_status( reg_status ),

    . reg_sa_p_clk_count_precharge( reg_sa_p_clk_count_precharge),

    . reg_sa_p_seq_n( reg_sa_p_seq_n),
    . reg_sa_p_seq0( reg_sa_p_seq0),
    . reg_sa_p_seq1( reg_sa_p_seq1),
    . reg_sa_p_seq2( reg_sa_p_seq2),
    . reg_sa_p_seq3( reg_sa_p_seq3),


    // outputs - sample acquisition
    . reg_adc_p_clk_count_aperture( reg_adc_p_clk_count_aperture),

    . reg_adc_p_clk_count_reset( reg_adc_p_clk_count_reset ),



/*


    .reg_adc_p_clk_count_reset(reg_adc_p_clk_count_reset ),

    // outputs adc
    .reg_adc_clk_count_refmux_reset({{ 8 { 1'b0 } }, adc2_clk_count_refmux_reset_last }  ) ,
    .reg_adc_clk_count_refmux_neg(  adc2_clk_count_refmux_neg_last   ) ,
    .reg_adc_clk_count_refmux_pos(  adc2_clk_count_refmux_pos_last  ) ,
    .reg_adc_clk_count_refmux_rd(  { {8{ 1'b0 }}, adc2_clk_count_refmux_rd_last }  ),
    .reg_adc_clk_count_mux_sig(                   adc2_clk_count_mux_sig_last   ),

    // adc stats
    .reg_adc_stat_count_refmux_pos_up( { {8{ 1'b0 }},adc2_stat_count_refmux_pos_up_last } ),
    .reg_adc_stat_count_refmux_neg_up( { {8{ 1'b0 }},adc2_stat_count_refmux_neg_up_last }),
    .reg_adc_stat_count_cmpr_cross_up(  { {8{ 1'b0 }},adc2_stat_count_cmpr_cross_up_last} )
*/
  );



endmodule


